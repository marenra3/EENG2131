`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Dunwoody College of Technology
// Engineer: Enrique Maritnez
// 
// Create Date: 12/01/2021 01:26:34 PM
// Design Name: 
// Module Name: wave_generator
// Project Name: audio generator 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module audio(
    input clk,
    output [7:0] JB);
    
    reg [9:0] sample_index;
    wire temp;
    
    wave_generator wg(clk,sample_index,{JB,temp});
    
    reg [9:0] count = 0;
    
    always@(posedge clk)
        begin
            if (count == 1000)
                begin
                 count <= 0;
                 if (sample_index == 1023)
                    begin
                     sample_index <= 0;
                    end
                  else
                   begin
                    sample_index = sample_index + 1;
                   end
                 
                end
             else
                begin
                 count <= count + 1;
                end
        end
endmodule
module audio_tb;
    reg clk = 0;
    wire [7:0] JB;
    
    integer i;
    
    audio test(clk,JB);
    
     initial begin
        for (i = 0; i <10000; i = i + 1)
        begin
        clk = ~clk;
        #10;
        end
    end
endmodule
    
module wave_generator(
    input clk,
    input [9:0] sample_index,
    output reg [8:0] sample = 0
    );
    reg [9:0] sine [0:1023];
    
    always@(posedge clk)
        begin
            sample<=sine[sample_index];
            
        end
    
     
    initial begin
    //case
        //0:8h'01;
        //
        sine[0] = 1;
        sine[1] = 3;
        sine[2] = 5;
        sine[3] = 7;
        sine[4] = 9;
        sine[5] = 11;
        sine[6] = 13;
        sine[7] = 15;
        sine[8] = 17;
        sine[9] = 19;
        sine[10] = 21;
        sine[11] = 23;
        sine[12] = 25;
        sine[13] = 27;
        sine[14] = 29;
        sine[15] = 31;
        sine[16] = 33;
        sine[17] = 35;
        sine[18] = 37;
        sine[19] = 39;
        sine[20] = 41;
        sine[21] = 43;
        sine[22] = 45;
        sine[23] = 47;
        sine[24] = 49;
        sine[25] = 51;
        sine[26] = 53;
        sine[27] = 55;
        sine[28] = 57;
        sine[29] = 59;
        sine[30] = 61;
        sine[31] = 63;
        sine[32] = 65;
        sine[33] = 67;
        sine[34] = 69;
        sine[35] = 71;
        sine[36] = 73;
        sine[37] = 75;
        sine[38]=77;
        sine[39]=79;
        sine[40]=81;
        sine[41]=83;
        sine[42]=85;
        sine[43]=87;
        sine[44]=89;
        sine[45]=91;
        sine[46]=93;
sine[47]=95;
sine[48]=97;
sine[49]=99;
sine[50]=101;
sine[51]=103;
sine[52]=105;
sine[53]=107;
sine[54]=109;
sine[55]=111;
sine[56]=113;
sine[57]=115;
sine[58]=117;
sine[59]=119;
sine[60]=121;
sine[61]=123;
sine[62]=125;
sine[63]=127;
sine[64]=129;
sine[65]=131;
sine[66]=133;
sine[67]=135;
sine[68]=137;
sine[69]=139;
sine[70]=141;
sine[71]=143;
sine[72]=145;
sine[73]=147;
sine[74]=149;
sine[75]=151;
sine[76]=153;
sine[77]=155;
sine[78]=157;
sine[79]=159;
sine[80]=161;
sine[81]=163;
sine[82]=165;
sine[83]=167;
sine[84]=169;
sine[85]=171;
sine[86]=173;
sine[87]=175;
sine[88]=177;
sine[89]=179;
sine[90]=181;
sine[91]=183;
sine[92]=185;
sine[93]=187;
sine[94]=189;
sine[95]=191;
sine[96]=193;
sine[97]=195;
sine[98]=197;
sine[99]=199;
sine[100]=201;
sine[101]=203;
sine[102]=205;
sine[103]=207;
sine[104]=209;
sine[105]=211;
sine[106]=213;
sine[107]=215;
sine[108]=217;
sine[109]=219;
sine[110]=221;
sine[111]=223;
sine[112]=225;
sine[113]=227;
sine[114]=229;
sine[115]=231;
sine[116]=233;
sine[117]=235;
sine[118]=237;
sine[119]=239;
sine[120]=241;
sine[121]=243;
sine[122]=245;
sine[123]=247;
sine[124]=249;
sine[125]=251;
sine[126]=253;
sine[127]=255;
sine[128]=257;
sine[129]=259;
sine[130]=261;
sine[131]=263;
sine[132]=265;
sine[133]=267;
sine[134]=269;
sine[135]=271;
sine[136]=273;
sine[137]=275;
sine[138]=277;
sine[139]=279;
sine[140]=281;
sine[141]=283;
sine[142]=285;
sine[143]=287;
sine[144]=289;
sine[145]=291;
sine[146]=293;
sine[147]=295;
sine[148] = 297;
sine[149] = 299;
sine[150] = 301;
sine[151] =303;
sine[152] = 305;
sine[153] = 307;
sine[154] = 309;
sine[155] = 311;
sine[156] = 313;
sine[157] = 315;
sine[158] = 317;
sine[159] = 319;
sine[160] = 321;
sine[161] = 323;
sine[162] = 325;
sine[163] = 327;
sine[164] = 329;
sine[165] = 331;
sine[166] = 333;	
sine [167]	=	335	;
sine [168]	=	337	;
sine [169]	=	339	;
sine [170]	=	341	;
sine [171]	=	343	;
sine [172]	=	345	;
sine [173]	=	347	;
sine [174]	=	349	;
sine [175]	=	351	;
sine [176]	=	353	;
sine [177]	=	355	;
sine [178]	=	357	;
sine [179]	=	359	;
sine [180]	=	361	;
sine [181]	=	363	;
sine [182]	=	365	;
sine [183]	=	367	;
sine [184]	=	369	;
sine [185]	=	371	;
sine [186]	=	373	;
sine [187]	=	375	;
sine [188]	=	377	;
sine [189]	=	379	;
sine [190]	=	381	;
sine [191]=	383	;
sine [192]=	385	;
sine [193]	=	387	;
sine [194]	=	389	;
sine [195]	=	391	;
sine [196]	=	393	;
sine [197]	=	395	;
sine [198]	=	397	;
sine [199]	=	399	;
sine [200]	=	401	;
sine [201]	=	403	;
sine [202]	=	405	;
sine [203]	=	407	;
sine [204]	=	409	;
sine [205]	=	411	;
sine [206]	=	413	;
sine [207]=	415	;
sine[208]=	417	;
sine [209]=	419	;
sine [210]=	421	;
sine [211]=	423	;
sine [212]	=	425	;
sine [213]	=	427	;
sine [214]	=	429	;
sine [215]	=	431	;
sine [216]	=	433	;
sine [217]	=	435	;
sine [218]	=	437	;
sine [219]	=	439	;
sine [220]	=	441	;
sine [221]	=	443	;
sine [222]	=	445	;
sine [223]	=	447	;
sine [224]	=	449	;
sine [225]	=	451	;
sine [226]	=	453	;
sine [227]	=	455	;
sine [228]	=	457	;
sine [229]	=	459	;
sine [230]=	461	;
sine	[	231	]	=	463	;
sine	[	232	]	=	465	;
sine	[	233	]	=	467	;
sine	[	234	]	=	469	;
sine	[	235	]	=	471	;
sine	[	236	]	=	473	;
sine	[	237	]	=	475	;
sine	[	238	]	=	477	;
sine	[	239	]	=	479	;
sine	[	240	]	=	481	;
sine	[	241	]	=	483	;
sine	[	242	]	=	485	;
sine	[	243	]	=	487	;
sine	[	244	]	=	489	;
sine	[	245	]	=	491	;
sine	[	246	]	=	493	;
sine	[	247	]	=	495	;
sine	[	248	]	=	497	;
sine	[	249	]	=	499	;
sine	[	250	]	=	501	;
sine	[	251	]	=	503	;
sine	[	252	]	=	505	;
sine	[	253	]	=	507	;
sine	[	254	]	=	509	;
sine	[	255	]	=	511	;
sine	[	256	]	=	513	;
sine	[	257	]	=	513	;
sine	[	258	]	=	511	;
sine	[	259	]	=	509	;
sine	[	260	]	=	507	;
sine	[	261	]	=	505	;
sine	[	262	]	=	503	;
sine	[	263	]	=	501	;
sine	[	264	]	=	499	;
sine	[	265	]	=	497	;
sine	[	266	]	=	495	;
sine	[	267	]	=	493	;
sine	[	268	]	=	491	;
sine	[	269	]	=	489	;
sine	[	270	]	=	487	;
sine	[	271	]	=	485	;
sine	[	272	]	=	483	;
sine	[	273	]	=	481	;
sine	[	274	]	=	479	;
sine	[	275	]	=	477	;
sine	[	276	]	=	475	;
sine	[	277	]	=	473	;
sine	[	278	]	=	471	;
sine	[	279	]	=	469	;
sine	[	280	]	=	467	;
sine	[	281	]	=	465	;
sine	[	282	]	=	463	;
sine	[	283	]	=	461	;
sine	[	284	]	=	459	;
sine	[	285	]	=	457	;
sine	[	286	]	=	455	;
sine	[	287	]	=	453	;
sine	[	288	]	=	451	;
sine	[	289	]	=	449	;
sine	[	290	]	=	447	;
sine	[	291	]	=	445	;
sine	[	292	]	=	443	;
sine	[	293	]	=	441	;
sine	[	294	]	=	439	;
sine	[	295	]	=	437	;
sine	[	296	]	=	435	;
sine	[	297	]	=	433	;
sine	[	298	]	=	431	;
sine	[	299	]	=	429	;
sine	[	300	]	=	427	;
sine	[	301	]	=	425	;
sine	[	302	]	=	423	;
sine	[	303	]	=	421	;
sine	[	304	]	=	419	;
sine	[	305	]	=	417	;
sine	[	306	]	=	415	;
sine	[	307	]	=	413	;
sine	[	308	]	=	411	;
sine	[	309	]	=	409	;
sine	[	310	]	=	407	;
sine	[	311	]	=	405	;
sine	[	312	]	=	403	;
sine	[	313	]	=	401	;
sine	[	314	]	=	399	;
sine	[	315	]	=	397	;
sine	[	316	]	=	395	;
sine	[	317	]	=	393	;
sine	[	318	]	=	391	;
sine	[	319	]	=	389	;
sine	[	320	]	=	387	;
sine	[	321	]	=	385	;
sine	[	322	]	=	383	;
sine	[	323	]	=	381	;
sine	[	324	]	=	379	;
sine	[	325	]	=	377	;
sine	[	326	]	=	375	;
sine	[	327	]	=	373	;
sine	[	328	]	=	371	;
sine	[	329	]	=	369	;
sine	[	330	]	=	367	;
sine	[	331	]	=	365	;
sine	[	332	]	=	363	;
sine	[	333	]	=	361	;
sine	[	334	]	=	359	;
sine	[	335	]	=	357	;
sine	[	336	]	=	355	;
sine	[	337	]	=	353	;
sine	[	338	]	=	351	;
sine	[	339	]	=	349	;
sine	[	340	]	=	347	;
sine	[	341	]	=	345	;
sine	[	342	]	=	343	;
sine	[	343	]	=	341	;
sine	[	344	]	=	339	;
sine	[	345	]	=	337	;
sine	[	346	]	=	335	;
sine	[	347	]	=	333	;
sine	[	348	]	=	331	;
sine	[	349	]	=	329	;
sine	[	350	]	=	327	;
sine	[	351	]	=	325	;
sine	[	352	]	=	323	;
sine	[	353	]	=	321	;
sine	[	354	]	=	319	;
sine	[	355	]	=	317	;
sine	[	356	]	=	315	;
sine	[	357	]	=	313	;
sine	[	358	]	=	311	;
sine	[	359	]	=	309	;
sine	[	360	]	=	307	;
sine	[	361	]	=	305	;
sine	[	362	]	=	303	;
sine	[	363	]	=	301	;
sine	[	364	]	=	299	;
sine	[	365	]	=	297	;
sine	[	366	]	=	295	;
sine	[	367	]	=	293	;
sine	[	368	]	=	291	;
sine	[	369	]	=	289	;
sine	[	370	]	=	287	;
sine	[	371	]	=	285	;
sine	[	372	]	=	283	;
sine	[	373	]	=	281	;
sine	[	374	]	=	279	;
sine	[	375	]	=	277	;
sine	[	376	]	=	275	;
sine	[	377	]	=	273	;
sine	[	378	]	=	271	;
sine	[	379	]	=	269	;
sine	[	380	]	=	267	;
sine	[	381	]	=	265	;
sine	[	382	]	=	263	;
sine	[	383	]	=	261	;
sine	[	384	]	=	259	;
sine	[	385	]	=	257	;
sine	[	386	]	=	255	;
sine	[	387	]	=	253	;
sine	[	388	]	=	251	;
sine	[	389	]	=	249	;
sine	[	390	]	=	247	;
sine	[	391	]	=	245	;
sine	[	392	]	=	243	;
sine	[	393	]	=	241	;
sine	[	394	]	=	239	;
sine	[	395	]	=	237	;
sine	[	396	]	=	235	;
sine	[	397	]	=	233	;
sine	[	398	]	=	231	;
sine	[	399	]	=	229	;
sine	[	400	]	=	227	;
sine	[	401	]	=	225	;
sine	[	402	]	=	223	;
sine	[	403	]	=	221	;
sine	[	404	]	=	219	;
sine	[	405	]	=	217	;
sine	[	406	]	=	215	;
sine	[	407	]	=	213	;
sine	[	408	]	=	211	;
sine	[	409	]	=	209	;
sine	[	410	]	=	207	;
sine	[	411	]	=	205	;
sine	[	412	]	=	203	;
sine	[	413	]	=	201	;
sine	[	414	]	=	199	;
sine	[	415	]	=	197	;
sine	[	416	]	=	195	;
sine	[	417	]	=	193	;
sine	[	418	]	=	191	;
sine	[	419	]	=	189	;
sine	[	420	]	=	187	;
sine	[	421	]	=	185	;
sine	[	422	]	=	183	;
sine	[	423	]	=	181	;
sine	[	424	]	=	179	;
sine	[	425	]	=	177	;
sine	[	426	]	=	175	;
sine	[	427	]	=	173	;
sine	[	428	]	=	171	;
sine	[	429	]	=	169	;
sine	[	430	]	=	167	;
sine	[	431	]	=	165	;
sine	[	432	]	=	163	;
sine	[	433	]	=	161	;
sine	[	434	]	=	159	;
sine	[	435	]	=	157	;
sine	[	436	]	=	155	;
sine	[	437	]	=	153	;
sine	[	438	]	=	151	;
sine	[	439	]	=	149	;
sine	[	440	]	=	147	;
sine	[	441	]	=	145	;
sine	[	442	]	=	143	;
sine	[	443	]	=	141	;
sine	[	444	]	=	139	;
sine	[	445	]	=	137	;
sine	[	446	]	=	135	;
sine	[	447	]	=	133	;
sine	[	448	]	=	131	;
sine	[	449	]	=	129	;
sine	[	450	]	=	127	;
sine	[	451	]	=	125	;
sine	[	452	]	=	123	;
sine	[	453	]	=	121	;
sine	[	454	]	=	119	;
sine	[	455	]	=	117	;
sine	[	456	]	=	115	;
sine	[	457	]	=	113	;
sine	[	458	]	=	111	;
sine	[	459	]	=	109	;
sine	[	460	]	=	107	;
sine	[	461	]	=	105	;
sine	[	462	]	=	103	;
sine	[	463	]	=	101	;
sine	[	464	]	=	99	;
sine	[	465	]	=	97	;
sine	[	466	]	=	95	;
sine	[	467	]	=	93	;
sine	[	468	]	=	91	;
sine	[	469	]	=	89	;
sine	[	470	]	=	87	;
sine	[	471	]	=	85	;
sine	[	472	]	=	83	;
sine	[	473	]	=	81	;
sine	[	474	]	=	79	;
sine	[	475	]	=	77	;
sine	[	476	]	=	75	;
sine	[	477	]	=	73	;
sine	[	478	]	=	71	;
sine	[	479	]	=	69	;
sine	[	480	]	=	67	;
sine	[	481	]	=	65	;
sine	[	482	]	=	63	;
sine	[	483	]	=	61	;
sine	[	484	]	=	59	;
sine	[	485	]	=	57	;
sine	[	486	]	=	55	;
sine	[	487	]	=	53	;
sine	[	488	]	=	51	;
sine	[	489	]	=	49	;
sine	[	490	]	=	47	;
sine	[	491	]	=	45	;
sine	[	492	]	=	43	;
sine	[	493	]	=	41	;
sine	[	494	]	=	39	;
sine	[	495	]	=	37	;
sine	[	496	]	=	35	;
sine	[	497	]	=	33	;
sine	[	498	]	=	31	;
sine	[	499	]	=	29	;
sine	[	500	]	=	27	;
sine	[	501	]	=	25	;
sine	[	502	]	=	23	;
sine	[	503	]	=	21	;
sine	[	504	]	=	19	;
sine	[	505	]	=	17	;
sine	[	506	]	=	15	;
sine	[	507	]	=	13	;
sine	[	508	]	=	11	;
sine	[	509	]	=	9	;
sine	[	510	]	=	7	;
sine	[	511	]	=	5	;
sine	[	512	]	=	3	;
sine	[	513	]	=	1	;
sine	[	514	]	=	-1	;
sine	[	515	]	=	-3	;
sine	[	516	]	=	-5	;
sine	[	517	]	=	-7	;
sine	[	518	]	=	-9	;
sine	[	519	]	=	-11	;
sine	[	520	]	=	-13	;
sine	[	521	]	=	-15	;
sine	[	522	]	=	-17	;
sine	[	523	]	=	-19	;
sine	[	524	]	=	-21	;
sine	[	525	]	=	-23	;
sine	[	526	]	=	-25	;
sine	[	527	]	=	-27	;
sine	[	528	]	=	-29	;
sine	[	529	]	=	-31	;
sine	[	530	]	=	-33	;
sine	[	531	]	=	-35	;
sine	[	532	]	=	-37	;
sine	[	533	]	=	-39	;
sine	[	534	]	=	-41	;
sine	[	535	]	=	-43	;
sine	[	536	]	=	-45	;
sine	[	537	]	=	-47	;
sine	[	538	]	=	-49	;
sine	[	539	]	=	-51	;
sine	[	540	]	=	-53	;
sine	[	541	]	=	-55	;
sine	[	542	]	=	-57	;
sine	[	543	]	=	-59	;
sine	[	544	]	=	-61	;
sine	[	545	]	=	-63	;
sine	[	546	]	=	-65	;
sine	[	547	]	=	-67	;
sine	[	548	]	=	-69	;
sine	[	549	]	=	-71	;
sine	[	550	]	=	-73	;
sine	[	551	]	=	-75	;
sine	[	552	]	=	-77	;
sine	[	553	]	=	-79	;
sine	[	554	]	=	-81	;
sine	[	555	]	=	-83	;
sine	[	556	]	=	-85	;
sine	[	557	]	=	-87	;
sine	[	558	]	=	-89	;
sine	[	559	]	=	-91	;
sine	[	560	]	=	-93	;
sine	[	561	]	=	-95	;
sine	[	562	]	=	-97	;
sine	[	563	]	=	-99	;
sine	[	564	]	=	-101	;
sine	[	565	]	=	-103	;
sine	[	566	]	=	-105	;
sine	[	567	]	=	-107	;
sine	[	568	]	=	-109	;
sine	[	569	]	=	-111	;
sine	[	570	]	=	-113	;
sine	[	571	]	=	-115	;
sine	[	572	]	=	-117	;
sine	[	573	]	=	-119	;
sine	[	574	]	=	-121	;
sine	[	575	]	=	-123	;
sine	[	576	]	=	-125	;
sine	[	577	]	=	-127	;
sine	[	578	]	=	-129	;
sine	[	579	]	=	-131	;
sine	[	580	]	=	-133	;
sine	[	581	]	=	-135	;
sine	[	582	]	=	-137	;
sine	[	583	]	=	-139	;
sine	[	584	]	=	-141	;
sine	[	585	]	=	-143	;
sine	[	586	]	=	-145	;
sine	[	587	]	=	-147	;
sine	[	588	]	=	-149	;
sine	[	589	]	=	-151	;
sine	[	590	]	=	-153	;
sine	[	591	]	=	-155	;
sine	[	592	]	=	-157	;
sine	[	593	]	=	-159	;
sine	[	594	]	=	-161	;
sine	[	595	]	=	-163	;
sine	[	596	]	=	-165	;
sine	[	597	]	=	-167	;
sine	[	598	]	=	-169	;
sine	[	599	]	=	-171	;
sine	[	600	]	=	-173	;
sine	[	601	]	=	-175	;
sine	[	602	]	=	-177	;
sine	[	603	]	=	-179	;
sine	[	604	]	=	-181	;
sine	[	605	]	=	-183	;
sine	[	606	]	=	-185	;
sine	[	607	]	=	-187	;
sine	[	608	]	=	-189	;
sine	[	609	]	=	-191	;
sine	[	610	]	=	-193	;
sine	[	611	]	=	-195	;
sine	[	612	]	=	-197	;
sine	[	613	]	=	-199	;
sine	[	614	]	=	-201	;
sine	[	615	]	=	-203	;
sine	[	616	]	=	-205	;
sine	[	617	]	=	-207	;
sine	[	618	]	=	-209	;
sine	[	619	]	=	-211	;
sine	[	620	]	=	-213	;
sine	[	621	]	=	-215	;
sine	[	622	]	=	-217	;
sine	[	623	]	=	-219	;
sine	[	624	]	=	-221	;
sine	[	625	]	=	-223	;
sine	[	626	]	=	-225	;
sine	[	627	]	=	-227	;
sine	[	628	]	=	-229	;
sine	[	629	]	=	-231	;
sine	[	630	]	=	-233	;
sine	[	631	]	=	-235	;
sine	[	632	]	=	-237	;
sine	[	633	]	=	-239	;
sine	[	634	]	=	-241	;
sine	[	635	]	=	-243	;
sine	[	636	]	=	-245	;
sine	[	637	]	=	-247	;
sine	[	638	]	=	-249	;
sine	[	639	]	=	-251	;
sine	[	640	]	=	-253	;
sine	[	641	]	=	-255	;
sine	[	642	]	=	-257	;
sine	[	643	]	=	-259	;
sine	[	644	]	=	-261	;
sine	[	645	]	=	-263	;
sine	[	646	]	=	-265	;
sine	[	647	]	=	-267	;
sine	[	648	]	=	-269	;
sine	[	649	]	=	-271	;
sine	[	650	]	=	-273	;
sine	[	651	]	=	-275	;
sine	[	652	]	=	-277	;
sine	[	653	]	=	-279	;
sine	[	654	]	=	-281	;
sine	[	655	]	=	-283	;
sine	[	656	]	=	-285	;
sine	[	657	]	=	-287	;
sine	[	658	]	=	-289	;
sine	[	659	]	=	-291	;
sine	[	660	]	=	-293	;
sine	[	661	]	=	-295	;
sine	[	662	]	=	-297	;
sine	[	663	]	=	-299	;
sine	[	664	]	=	-301	;
sine	[	665	]	=	-303	;
sine	[	666	]	=	-305	;
sine	[	667	]	=	-307	;
sine	[	668	]	=	-309	;
sine	[	669	]	=	-311	;
sine	[	670	]	=	-313	;
sine	[	671	]	=	-315	;
sine	[	672	]	=	-317	;
sine	[	673	]	=	-319	;
sine	[	674	]	=	-321	;
sine	[	675	]	=	-323	;
sine	[	676	]	=	-325	;
sine	[	677	]	=	-327	;
sine	[	678	]	=	-329	;
sine	[	679	]	=	-331	;
sine	[	680	]	=	-333	;
sine	[	681	]	=	-335	;
sine	[	682	]	=	-337	;
sine	[	683	]	=	-339	;
sine	[	684	]	=	-341	;
sine	[	685	]	=	-343	;
sine	[	686	]	=	-345	;
sine	[	687	]	=	-347	;
sine	[	688	]	=	-349	;
sine	[	689	]	=	-351	;
sine	[	690	]	=	-353	;
sine	[	691	]	=	-355	;
sine	[	692	]	=	-357	;
sine	[	693	]	=	-359	;
sine	[	694	]	=	-361	;
sine	[	695	]	=	-363	;
sine	[	696	]	=	-365	;
sine	[	697	]	=	-367	;
sine	[	698	]	=	-369	;
sine	[	699	]	=	-371	;
sine	[	700	]	=	-373	;
sine	[	701	]	=	-375	;
sine	[	702	]	=	-377	;
sine	[	703	]	=	-379	;
sine	[	704	]	=	-381	;
sine	[	705	]	=	-383	;
sine	[	706	]	=	-385	;
sine	[	707	]	=	-387	;
sine	[	708	]	=	-389	;
sine	[	709	]	=	-391	;
sine	[	710	]	=	-393	;
sine	[	711	]	=	-395	;
sine	[	712	]	=	-397	;
sine	[	713	]	=	-399	;
sine	[	714	]	=	-401	;
sine	[	715	]	=	-403	;
sine	[	716	]	=	-405	;
sine	[	717	]	=	-407	;
sine	[	718	]	=	-409	;
sine	[	719	]	=	-411	;
sine	[	720	]	=	-413	;
sine	[	721	]	=	-415	;
sine	[	722	]	=	-417	;
sine	[	723	]	=	-419	;
sine	[	724	]	=	-421	;
sine	[	725	]	=	-423	;
sine	[	726	]	=	-425	;
sine	[	727	]	=	-427	;
sine	[	728	]	=	-429	;
sine	[	729	]	=	-431	;
sine	[	730	]	=	-433	;
sine	[	731	]	=	-435	;
sine	[	732	]	=	-437	;
sine	[	733	]	=	-439	;
sine	[	734	]	=	-441	;
sine	[	735	]	=	-443	;
sine	[	736	]	=	-445	;
sine	[	737	]	=	-447	;
sine	[	738	]	=	-449	;
sine	[	739	]	=	-451	;
sine	[	740	]	=	-453	;
sine	[	741	]	=	-455	;
sine	[	742	]	=	-457	;
sine	[	743	]	=	-459	;
sine	[	744	]	=	-461	;
sine	[	745	]	=	-463	;
sine	[	746	]	=	-465	;
sine	[	747	]	=	-467	;
sine	[	748	]	=	-469	;
sine	[	749	]	=	-471	;
sine	[	750	]	=	-473	;
sine	[	751	]	=	-475	;
sine	[	752	]	=	-477	;
sine	[	753	]	=	-479	;
sine	[	754	]	=	-481	;
sine	[	755	]	=	-483	;
sine	[	756	]	=	-485	;
sine	[	757	]	=	-487	;
sine	[	758	]	=	-489	;
sine	[	759	]	=	-491	;
sine	[	760	]	=	-493	;
sine	[	761	]	=	-495	;
sine	[	762	]	=	-497	;
sine	[	763	]	=	-499	;
sine	[	764	]	=	-501	;
sine	[	765	]	=	-503	;
sine	[	766	]	=	-505	;
sine	[	767	]	=	-507	;
sine	[	768	]	=	-509	;
sine	[	769	]	=	-509	;
sine	[	770	]	=	-507	;
sine	[	771	]	=	-505	;
sine	[	772	]	=	-503	;
sine	[	773	]	=	-501	;
sine	[	774	]	=	-499	;
sine	[	775	]	=	-497	;
sine	[	776	]	=	-495	;
sine	[	777	]	=	-493	;
sine	[	778	]	=	-491	;
sine	[	779	]	=	-489	;
sine	[	780	]	=	-487	;
sine	[	781	]	=	-485	;
sine	[	782	]	=	-483	;
sine	[	783	]	=	-481	;
sine	[	784	]	=	-479	;
sine	[	785	]	=	-477	;
sine	[	786	]	=	-475	;
sine	[	787	]	=	-473	;
sine	[	788	]	=	-471	;
sine	[	789	]	=	-469	;
sine	[	790	]	=	-467	;
sine	[	791	]	=	-465	;
sine	[	792	]	=	-463	;
sine	[	793	]	=	-461	;
sine	[	794	]	=	-459	;
sine	[	795	]	=	-457	;
sine	[	796	]	=	-455	;
sine	[	797	]	=	-453	;
sine	[	798	]	=	-451	;
sine	[	799	]	=	-449	;
sine	[	800	]	=	-447	;
sine	[	801	]	=	-445	;
sine	[	802	]	=	-443	;
sine	[	803	]	=	-441	;
sine	[	804	]	=	-439	;
sine	[	805	]	=	-437	;
sine	[	806	]	=	-435	;
sine	[	807	]	=	-433	;
sine	[	808	]	=	-431	;
sine	[	809	]	=	-429	;
sine	[	810	]	=	-427	;
sine	[	811	]	=	-425	;
sine	[	812	]	=	-423	;
sine	[	813	]	=	-421	;
sine	[	814	]	=	-419	;
sine	[	815	]	=	-417	;
sine	[	816	]	=	-415	;
sine	[	817	]	=	-413	;
sine	[	818	]	=	-411	;
sine	[	819	]	=	-409	;
sine	[	820	]	=	-407	;
sine	[	821	]	=	-405	;
sine	[	822	]	=	-403	;
sine	[	823	]	=	-401	;
sine	[	824	]	=	-399	;
sine	[	825	]	=	-397	;
sine	[	826	]	=	-395	;
sine	[	827	]	=	-393	;
sine	[	828	]	=	-391	;
sine	[	829	]	=	-389	;
sine	[	830	]	=	-387	;
sine	[	831	]	=	-385	;
sine	[	832	]	=	-383	;
sine	[	833	]	=	-381	;
sine	[	834	]	=	-379	;
sine	[	835	]	=	-377	;
sine	[	836	]	=	-375	;
sine	[	837	]	=	-373	;
sine	[	838	]	=	-371	;
sine	[	839	]	=	-369	;
sine	[	840	]	=	-367	;
sine	[	841	]	=	-365	;
sine	[	842	]	=	-363	;
sine	[	843	]	=	-361	;
sine	[	844	]	=	-359	;
sine	[	845	]	=	-357	;
sine	[	846	]	=	-355	;
sine	[	847	]	=	-353	;
sine	[	848	]	=	-351	;
sine	[	849	]	=	-349	;
sine	[	850	]	=	-347	;
sine	[	851	]	=	-345	;
sine	[	852	]	=	-343	;
sine	[	853	]	=	-341	;
sine	[	854	]	=	-339	;
sine	[	855	]	=	-337	;
sine	[	856	]	=	-335	;
sine	[	857	]	=	-333	;
sine	[	858	]	=	-331	;
sine	[	859	]	=	-329	;
sine	[	860	]	=	-327	;
sine	[	861	]	=	-325	;
sine	[	862	]	=	-323	;
sine	[	863	]	=	-321	;
sine	[	864	]	=	-319	;
sine	[	865	]	=	-317	;
sine	[	866	]	=	-315	;
sine	[	867	]	=	-313	;
sine	[	868	]	=	-311	;
sine	[	869	]	=	-309	;
sine	[	870	]	=	-307	;
sine	[	871	]	=	-305	;
sine	[	872	]	=	-303	;
sine	[	873	]	=	-301	;
sine	[	874	]	=	-299	;
sine	[	875	]	=	-297	;
sine	[	876	]	=	-295	;
sine	[	877	]	=	-293	;
sine	[	878	]	=	-291	;
sine	[	879	]	=	-289	;
sine	[	880	]	=	-287	;
sine	[	881	]	=	-285	;
sine	[	882	]	=	-283	;
sine	[	883	]	=	-281	;
sine	[	884	]	=	-279	;
sine	[	885	]	=	-277	;
sine	[	886	]	=	-275	;
sine	[	887	]	=	-273	;
sine	[	888	]	=	-271	;
sine	[	889	]	=	-269	;
sine	[	890	]	=	-267	;
sine	[	891	]	=	-265	;
sine	[	892	]	=	-263	;
sine	[	893	]	=	-261	;
sine	[	894	]	=	-259	;
sine	[	895	]	=	-257	;
sine	[	896	]	=	-255	;
sine	[	897	]	=	-253	;
sine	[	898	]	=	-251	;
sine	[	899	]	=	-249	;
sine	[	900	]	=	-247	;
sine	[	901	]	=	-245	;
sine	[	902	]	=	-243	;
sine	[	903	]	=	-241	;
sine	[	904	]	=	-239	;
sine	[	905	]	=	-237	;
sine	[	906	]	=	-235	;
sine	[	907	]	=	-233	;
sine	[	908	]	=	-231	;
sine	[	909	]	=	-229	;
sine	[	910	]	=	-227	;
sine	[	911	]	=	-225	;
sine	[	912	]	=	-223	;
sine	[	913	]	=	-221	;
sine	[	914	]	=	-219	;
sine	[	915	]	=	-217	;
sine	[	916	]	=	-215	;
sine	[	917	]	=	-213	;
sine	[	918	]	=	-211	;
sine	[	919	]	=	-209	;
sine	[	920	]	=	-207	;
sine	[	921	]	=	-205	;
sine	[	922	]	=	-203	;
sine	[	923	]	=	-201	;
sine	[	924	]	=	-199	;
sine	[	925	]	=	-197	;
sine	[	926	]	=	-195	;
sine	[	927	]	=	-193	;
sine	[	928	]	=	-191	;
sine	[	929	]	=	-189	;
sine	[	930	]	=	-187	;
sine	[	931	]	=	-185	;
sine	[	932	]	=	-183	;
sine	[	933	]	=	-181	;
sine	[	934	]	=	-179	;
sine	[	935	]	=	-177	;
sine	[	936	]	=	-175	;
sine	[	937	]	=	-173	;
sine	[	938	]	=	-171	;
sine	[	939	]	=	-169	;
sine	[	940	]	=	-167	;
sine	[	941	]	=	-165	;
sine	[	942	]	=	-163	;
sine	[	943	]	=	-161	;
sine	[	944	]	=	-159	;
sine	[	945	]	=	-157	;
sine	[	946	]	=	-155	;
sine	[	947	]	=	-153	;
sine	[	948	]	=	-151	;
sine	[	949	]	=	-149	;
sine	[	950	]	=	-147	;
sine	[	951	]	=	-145	;
sine	[	952	]	=	-143	;
sine	[	953	]	=	-141	;
sine	[	954	]	=	-139	;
sine	[	955	]	=	-137	;
sine	[	956	]	=	-135	;
sine	[	957	]	=	-133	;
sine	[	958	]	=	-131	;
sine	[	959	]	=	-129	;
sine	[	960	]	=	-127	;
sine	[	961	]	=	-125	;
sine	[	962	]	=	-123	;
sine	[	963	]	=	-121	;
sine	[	964	]	=	-119	;
sine	[	965	]	=	-117	;
sine	[	966	]	=	-115	;
sine	[	967	]	=	-113	;
sine	[	968	]	=	-111	;
sine	[	969	]	=	-109	;
sine	[	970	]	=	-107	;
sine	[	971	]	=	-105	;
sine	[	972	]	=	-103	;
sine	[	973	]	=	-101	;
sine	[	974	]	=	-99	;
sine	[	975	]	=	-97	;
sine	[	976	]	=	-95	;
sine	[	977	]	=	-93	;
sine	[	978	]	=	-91	;
sine	[	979	]	=	-89	;
sine	[	980	]	=	-87	;
sine	[	981	]	=	-85	;
sine	[	982	]	=	-83	;
sine	[	983	]	=	-81	;
sine	[	984	]	=	-79	;
sine	[	985	]	=	-77	;
sine	[	986	]	=	-75	;
sine	[	987	]	=	-73	;
sine	[	988	]	=	-71	;
sine	[	989	]	=	-69	;
sine	[	990	]	=	-67	;
sine	[	991	]	=	-65	;
sine	[	992	]	=	-63	;
sine	[	993	]	=	-61	;
sine	[	994	]	=	-59	;
sine	[	995	]	=	-57	;
sine	[	996	]	=	-55	;
sine	[	997	]	=	-53	;
sine	[	998	]	=	-51	;
sine	[	999	]	=	-49	;
sine	[	1000	]	=	-47	;
sine	[	1001	]	=	-45	;
sine	[	1002	]	=	-43	;
sine	[	1003	]	=	-41	;
sine	[	1004	]	=	-39	;
sine	[	1005	]	=	-37	;
sine	[	1006	]	=	-35	;
sine	[	1007	]	=	-33	;
sine	[	1008	]	=	-31	;
sine	[	1009	]	=	-29	;
sine	[	1010	]	=	-27	;
sine	[	1011	]	=	-25	;
sine	[	1012	]	=	-23	;
sine	[	1013	]	=	-21	;
sine	[	1014	]	=	-19	;
sine	[	1015	]	=	-17	;
sine	[	1016	]	=	-15	;
sine	[	1017	]	=	-13	;
sine	[	1018	]	=	-11	;
sine	[	1019	]	=	-9	;
sine	[	1020	]	=	-7	;
sine	[	1021	]	=	-5	;
sine	[	1022	]	=	-3	;
sine	[	1023	]	=	-1	;



end
//if (counter == sw) begin
//            JB <= JB + 1;
//            counter <= 0;
//        end else begin
//            counter <= counter + 1;

endmodule
//module wave_generator_tb;
//    reg clk;
//    reg [9:0] sample_index;
//    wire [8:0] sample;
    
    
//    wave_generator dut(clk,sample_index,sample);
    
     
//     initial begin
       
        
//        sample_index = 9'b000000011;
//        #10;
//        sample_index = 9'b000011001;
//        #10;
//        sample_index = 9'b000101010; 
//        #10;
//        sample_index = 9'b001101001; 
//        #10;
//        sample_index = 9'b001101110; 
//        #10;
//        sample_index = 9'b010000010; 
//        #10;
//        sample_index = 9'b011101010; 
//        #10;
//        sample_index = 9'b100101101;
//        #10; 
        
//    end
//endmodule  
//module accumod (in, acc, clk, reset);

//input [7:0] in;

//input clk, reset;

//output [7:0] acc;

//reg [7:0] acc;

//always@(clk) begin

//if(reset)

//acc <= 8'b00000000;

//else

//acc <= acc + in;

//end

//endmodule 
// input clk,
//    output reg [7:0] JB
//    );
    
//    reg [7:0] sine [0:29];
//    integer i;  
//     always @(posedge(clk))
//    begin
//        JB = sine[i];
//        i <= i+ 1;

//module wave_generator_tb;
//   reg clk;
//   wire [7:0] JB;

//   wave_generator test(clk,JB);

//   initial clk = 0;
//   always #10 clk = ~clk;
    
//endmodule